module(
input a,
input b,
input s,
input c
);
assign c=s?a:b;
endmodule
