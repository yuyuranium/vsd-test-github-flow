module test;
   
endmodule
