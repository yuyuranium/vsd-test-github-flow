module test;

endmodule
